module flip_flop_d(
	input d,
	output q, nq
);



endmodule