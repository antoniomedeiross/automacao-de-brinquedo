module debounce(
	input clk, pulso, 
	output signal
);	
// clock de 50 Hz
	wire fios_saidaff1;

	flip_flop_d ff1 ();
	flip_flop_d ff2 ();

endmodule